`timescale 1ns / 1ps
// Single Port ROM

module single_port_rom
#(parameter DATA_WIDTH=96, parameter ADDR_WIDTH=12)
(
	input [(ADDR_WIDTH-1):0] addr,
	input clk, 
	output reg [(DATA_WIDTH-1):0] q
);

	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

	initial
	begin
		$readmemb("single_port_rom_init.mem", rom);
	end

	always @ (posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
